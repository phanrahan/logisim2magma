module main (input [0:1] SWITCH, output [0:3] LED);
wire inst0_Q;
wire inst1_O;
wire inst2_Q;
wire inst3_O;
wire inst4_O;
wire inst5_O;
wire inst6_O;
wire inst7_Q;
wire inst8_O;
wire inst9_O;
wire inst10_O;
wire inst11_O;
wire inst12_O;
wire inst13_O;
wire inst14_Q;
wire inst15_O;
wire inst16_O;
wire inst17_O;
FDRSE #(.INIT(1'b0)) inst0 (.CE(1'b1), .R(1'b0), .S(1'b0), .D(inst1_O), .Q(inst0_Q));
LUT2 #(.INIT(4'h6)) inst1 (.I0(inst0_Q), .I1(inst12_O), .O(inst1_O));
FDRSE #(.INIT(1'b0)) inst2 (.CE(1'b1), .R(1'b0), .S(1'b0), .D(inst3_O), .Q(inst2_Q));
LUT2 #(.INIT(4'h6)) inst3 (.I0(inst2_Q), .I1(inst6_O), .O(inst3_O));
LUT2 #(.INIT(4'h8)) inst4 (.I0(inst13_O), .I1(inst0_Q), .O(inst4_O));
LUT2 #(.INIT(4'h8)) inst5 (.I0(inst4_O), .I1(inst7_Q), .O(inst5_O));
LUT2 #(.INIT(4'hE)) inst6 (.I0(inst5_O), .I1(inst16_O), .O(inst6_O));
FDRSE #(.INIT(1'b0)) inst7 (.CE(1'b1), .R(1'b0), .S(1'b0), .D(inst8_O), .Q(inst7_Q));
LUT2 #(.INIT(4'h6)) inst8 (.I0(inst7_Q), .I1(inst11_O), .O(inst8_O));
LUT1 #(.INIT(2'h1)) inst9 (.I0(SWITCH[0]), .O(inst9_O));
LUT2 #(.INIT(4'hF)) inst10 (.I0(inst14_Q), .I1(inst9_O), .O(inst10_O));
LUT2 #(.INIT(4'hE)) inst11 (.I0(inst4_O), .I1(inst17_O), .O(inst11_O));
LUT2 #(.INIT(4'hE)) inst12 (.I0(inst13_O), .I1(inst10_O), .O(inst12_O));
LUT2 #(.INIT(4'h8)) inst13 (.I0(SWITCH[0]), .I1(inst14_Q), .O(inst13_O));
FDRSE #(.INIT(1'b0)) inst14 (.CE(1'b1), .R(1'b0), .S(1'b0), .D(inst15_O), .Q(inst14_Q));
LUT2 #(.INIT(4'h6)) inst15 (.I0(inst14_Q), .I1(1'b1), .O(inst15_O));
LUT2 #(.INIT(4'hF)) inst16 (.I0(inst7_Q), .I1(inst17_O), .O(inst16_O));
LUT2 #(.INIT(4'hF)) inst17 (.I0(inst0_Q), .I1(inst10_O), .O(inst17_O));
assign LED = {inst14_Q, inst0_Q, inst7_Q, inst2_Q};
endmodule

